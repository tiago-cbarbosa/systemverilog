$ -> tasks
$dysplay("Hello, my value in decimal is %d", var_a)
$finish
$stop
$exit
$time - ex $display("Simulation error at time %t in output a with value %d", out_a);
$random